-- megafunction wizard: %ALTFP_EXP%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTFP_EXP 

-- ============================================================
-- File Name: f_p_exp.vhd
-- Megafunction Name(s):
-- 			ALTFP_EXP
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2018  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details.


--altfp_exp CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="MAX 10" PIPELINE=17 ROUNDING="TO_NEAREST" WIDTH_EXP=8 WIDTH_MAN=23 clock data result
--VERSION_BEGIN 18.1 cbx_altfp_exp 2018:09:12:13:04:09:SJ cbx_altmult_opt 2018:09:12:13:04:09:SJ cbx_cycloneii 2018:09:12:13:04:09:SJ cbx_lpm_add_sub 2018:09:12:13:04:09:SJ cbx_lpm_clshift 2018:09:12:13:04:09:SJ cbx_lpm_compare 2018:09:12:13:04:09:SJ cbx_lpm_mult 2018:09:12:13:04:09:SJ cbx_lpm_mux 2018:09:12:13:04:09:SJ cbx_mgl 2018:09:12:14:15:07:SJ cbx_nadder 2018:09:12:13:04:09:SJ cbx_padd 2018:09:12:13:04:09:SJ cbx_stratix 2018:09:12:13:04:09:SJ cbx_stratixii 2018:09:12:13:04:09:SJ cbx_util_mgl 2018:09:12:13:04:09:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.lpm_components.all;

--synthesis_resources = lpm_add_sub 9 lpm_clshift 1 lpm_compare 3 lpm_mult 5 lpm_mux 3 mux21 124 reg 745 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  f_p_exp_altfp_exp_jmc IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END f_p_exp_altfp_exp_jmc;

 ARCHITECTURE RTL OF f_p_exp_altfp_exp_jmc IS

	 SIGNAL	 barrel_shifter_underflow_dffe2_15_pipes0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_15_pipes1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_15_pipes2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_15_pipes3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_15_pipes4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_15_pipes5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_15_pipes6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_15_pipes7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_15_pipes8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_15_pipes9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_15_pipes10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_15_pipes11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_15_pipes12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_15_pipes13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 barrel_shifter_underflow_dffe2_15_pipes14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_15_pipes0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_15_pipes1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_15_pipes2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_15_pipes3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_15_pipes4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_15_pipes5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_15_pipes6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_15_pipes7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_15_pipes8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_15_pipes9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_15_pipes10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_15_pipes11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_15_pipes12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_15_pipes13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 distance_overflow_dffe2_15_pipes14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_0	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_1	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_10	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_2	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_3	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_4	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_5	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_6	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_7	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_8	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_b4_bias_dffe_9	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_value_dffe1	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 extra_ln2_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 extra_ln2_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 extra_ln2_dffe_2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 extra_ln2_dffe_3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 extra_ln2_dffe_4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 extra_ln2_dffe_5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_extra_ln2_dffe_5_w_lg_q157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 fraction_dffe1	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_16_pipes0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_16_pipes1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_16_pipes2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_16_pipes3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_16_pipes4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_16_pipes5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_16_pipes6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_16_pipes7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_16_pipes8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_16_pipes9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_16_pipes10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_16_pipes11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_16_pipes12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_16_pipes13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_16_pipes14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_16_pipes15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_16_pipes0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_16_pipes1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_16_pipes2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_16_pipes3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_16_pipes4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_16_pipes5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_16_pipes6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_16_pipes7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_16_pipes8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_16_pipes9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_16_pipes10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_16_pipes11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_16_pipes12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_16_pipes13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_16_pipes14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_16_pipes15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_16_pipes0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_16_pipes1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_16_pipes2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_16_pipes3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_16_pipes4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_16_pipes5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_16_pipes6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_16_pipes7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_16_pipes8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_16_pipes9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_16_pipes10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_16_pipes11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_16_pipes12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_16_pipes13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_16_pipes14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_16_pipes15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_overflow_dffe15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_prod_dffe14	:	STD_LOGIC_VECTOR(61 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_round_dffe15	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 result_pipe_dffe16	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 round_up_dffe15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_sign_dffe_w_lg_q448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_sign_dffe_w_lg_q434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 tbl1_compare_dffe11_4_pipes0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 tbl1_compare_dffe11_4_pipes1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 tbl1_compare_dffe11_4_pipes2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 tbl1_compare_dffe11_4_pipes3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 tbl1_tbl2_prod_dffe12	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 tbl3_taylor_prod_dffe12	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_fixed_dffe_0	:	STD_LOGIC_VECTOR(37 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_fixed_dffe_1	:	STD_LOGIC_VECTOR(37 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_fixed_dffe_2	:	STD_LOGIC_VECTOR(37 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_fixed_dffe_3	:	STD_LOGIC_VECTOR(37 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_fixed_dffe_4	:	STD_LOGIC_VECTOR(37 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 xf_pre_2_dffe10	:	STD_LOGIC_VECTOR(37 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 xf_pre_dffe9	:	STD_LOGIC_VECTOR(37 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 xi_exp_value_dffe4	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 xi_ln2_prod_dffe7	:	STD_LOGIC_VECTOR(45 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 xi_prod_dffe3	:	STD_LOGIC_VECTOR(20 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exp_minus_bias_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exp_minus_bias_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exp_minus_bias_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exp_value_add_bias_w_lg_w_result_range445w446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_value_add_bias_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exp_value_add_bias_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exp_value_add_bias_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exp_value_add_bias_w_result_range445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_value_man_over_w_lg_w_lg_w_result_range435w436w437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_value_man_over_w_lg_w_result_range435w436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_value_man_over_w_lg_w_lg_w_lg_w_result_range435w436w437w438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_value_man_over_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exp_value_man_over_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exp_value_man_over_w_result_range435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_invert_exp_value_dataa	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_invert_exp_value_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_invert_exp_value_w_result_range130w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_man_round_datab	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_man_round_result	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_one_minus_xf_dataa	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_one_minus_xf_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_x_fixed_minus_xiln2_datab	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_x_fixed_minus_xiln2_result	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_xf_minus_ln2_datab	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_xf_minus_ln2_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_xi_add_one_datab	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_xi_add_one_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_result	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_distance_overflow_comp_agb	:	STD_LOGIC;
	 SIGNAL  wire_tbl1_compare_ageb	:	STD_LOGIC;
	 SIGNAL  wire_underflow_compare_agb	:	STD_LOGIC;
	 SIGNAL  wire_man_prod_result	:	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  wire_tbl1_tbl2_prod_result	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_datab	:	STD_LOGIC_VECTOR (29 DOWNTO 0);
	 SIGNAL  wire_tbl3_taylor_prod_result	:	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  wire_xi_ln2_prod_result	:	STD_LOGIC_VECTOR (45 DOWNTO 0);
	 SIGNAL  wire_xi_prod_result	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_table_one_data_2d	:	STD_LOGIC_2D(31 DOWNTO 0, 31 DOWNTO 0);
	 SIGNAL  wire_table_one_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_table_three_data_2d	:	STD_LOGIC_2D(31 DOWNTO 0, 20 DOWNTO 0);
	 SIGNAL  wire_table_three_result	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_table_two_data_2d	:	STD_LOGIC_2D(31 DOWNTO 0, 25 DOWNTO 0);
	 SIGNAL  wire_table_two_result	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL	wire_cin_to_bias_dataout	:	STD_LOGIC;
	 SIGNAL	wire_exp_result_mux_prea_dataout	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL  wire_exp_result_mux_prea_w_lg_dataout557w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	wire_exp_value_b4_biasa_dataout	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	wire_exp_value_selecta_dataout	:	STD_LOGIC_VECTOR(5 DOWNTO 0);
	 SIGNAL	wire_exp_value_to_compare_muxa_dataout	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	wire_exp_value_to_ln2a_dataout	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	wire_extra_ln2_muxa_dataout	:	STD_LOGIC_VECTOR(30 DOWNTO 0);
	 SIGNAL	wire_man_result_muxa_dataout	:	STD_LOGIC_VECTOR(22 DOWNTO 0);
	 SIGNAL	wire_xf_muxa_dataout	:	STD_LOGIC_VECTOR(30 DOWNTO 0);
	 SIGNAL  wire_w_lg_man_prod_shifted408w	:	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  wire_w_lg_man_prod_wire407w	:	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  wire_w_lg_underflow_w554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range10w34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range13w36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range16w38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range19w40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range22w42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range25w44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range28w46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_data_all_one_w_range47w119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range563w564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range568w569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range573w574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range578w579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range583w584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range588w589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range593w594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range492w493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range495w496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range498w499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range501w502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range504w505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range507w508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range510w511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range513w514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range516w517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range519w520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range465w466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range522w523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range525w526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range528w529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range468w469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range471w472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range474w475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range477w478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range480w481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range483w484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range486w487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_round_wi_range489w490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_underflow_w554w555w556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_barrel_shifter_underflow553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_is_infinity_wo443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_is_nan_wo442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_is_zero_wo444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_underflow_w454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_data_not_zero_w_range116w118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_prod_wo_range402w406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_underflow_w554w555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w551w552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_overflow_w536w537w538w539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_overflow_w536w537w538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_barrel_shifter_underflow549w550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_overflow_w542w543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_overflow_w536w537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_barrel_shifter_underflow549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_distance_overflow447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_distance_overflow456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_overflow_w542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_overflow_w536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range78w79w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range81w82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range84w85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range87w88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range90w91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range93w94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range96w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range99w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range102w103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range105w106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range51w52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range108w109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range111w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range114w115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range10w11w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range13w14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range16w17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range19w20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range22w23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range25w26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range54w55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range28w29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range57w58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range60w61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range63w64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range66w67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range69w70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range72w73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_data_range75w76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range563w566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range568w571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range573w576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range578w581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range583w586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range588w591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_result_w_range593w595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_prod_result_range424w425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_prod_result_range421w422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_prod_result_range418w419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_prod_result_range415w416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  addr_val_more_than_one :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  barrel_shifter_data :	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  barrel_shifter_distance :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  barrel_shifter_underflow :	STD_LOGIC;
	 SIGNAL  barrel_shifter_underflow_wi :	STD_LOGIC;
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  distance_overflow :	STD_LOGIC;
	 SIGNAL  distance_overflow_val_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  distance_overflow_wi :	STD_LOGIC;
	 SIGNAL  exp_bias :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_bias_all_ones_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_data_all_one_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_data_not_zero_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_invert :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_one :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_out_all_one_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_out_not_zero_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_result_out :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_result_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_value :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_value_wi :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_value_wo :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  extra_ln2 :	STD_LOGIC;
	 SIGNAL  fraction :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  fraction_wi :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  fraction_wo :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  gnd_w :	STD_LOGIC;
	 SIGNAL  guard_bit :	STD_LOGIC;
	 SIGNAL  input_is_infinity_wi :	STD_LOGIC;
	 SIGNAL  input_is_infinity_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_wo :	STD_LOGIC;
	 SIGNAL  input_is_zero_wi :	STD_LOGIC;
	 SIGNAL  input_is_zero_wo :	STD_LOGIC;
	 SIGNAL  ln2_w :	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  man_data_not_zero_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_overflow :	STD_LOGIC;
	 SIGNAL  man_overflow_wi :	STD_LOGIC;
	 SIGNAL  man_overflow_wo :	STD_LOGIC;
	 SIGNAL  man_prod_result :	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  man_prod_shifted :	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  man_prod_wi :	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  man_prod_wire :	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  man_prod_wo :	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  man_result_all_ones :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_result_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_round_wi :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_round_wo :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  nan_w :	STD_LOGIC;
	 SIGNAL  negative_infinity :	STD_LOGIC;
	 SIGNAL  one_over_ln2_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  overflow_w :	STD_LOGIC;
	 SIGNAL  positive_infinity :	STD_LOGIC;
	 SIGNAL  result_pipe_wi :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  result_pipe_wo :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  result_underflow_w :	STD_LOGIC;
	 SIGNAL  round_bit :	STD_LOGIC;
	 SIGNAL  round_up :	STD_LOGIC;
	 SIGNAL  round_up_wi :	STD_LOGIC;
	 SIGNAL  round_up_wo :	STD_LOGIC;
	 SIGNAL  shifted_value :	STD_LOGIC;
	 SIGNAL  sign_w :	STD_LOGIC;
	 SIGNAL  sticky_bits :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  table_one_data :	STD_LOGIC_VECTOR (1023 DOWNTO 0);
	 SIGNAL  table_one_out :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  table_three_data :	STD_LOGIC_VECTOR (671 DOWNTO 0);
	 SIGNAL  table_three_out :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  table_three_out_tmp :	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  table_two_data :	STD_LOGIC_VECTOR (831 DOWNTO 0);
	 SIGNAL  table_two_out :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  table_two_out_tmp :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  tbl1_compare_wi :	STD_LOGIC;
	 SIGNAL  tbl1_compare_wo :	STD_LOGIC;
	 SIGNAL  tbl1_tbl2_prod_wi :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  tbl1_tbl2_prod_wo :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  tbl3_taylor_prod_wi :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  tbl3_taylor_prod_wo :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  underflow_compare_val_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  underflow_w :	STD_LOGIC;
	 SIGNAL  x_fixed :	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  xf :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  xf_pre :	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  xf_pre_2_wi :	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  xf_pre_2_wo :	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  xf_pre_wi :	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  xf_pre_wo :	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  xi_exp_value :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  xi_exp_value_wi :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  xi_exp_value_wo :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  xi_ln2_prod_wi :	STD_LOGIC_VECTOR (45 DOWNTO 0);
	 SIGNAL  xi_ln2_prod_wo :	STD_LOGIC_VECTOR (45 DOWNTO 0);
	 SIGNAL  xi_prod_wi :	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  xi_prod_wo :	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_w_data_range78w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range81w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range84w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range16w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_range75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_all_one_w_range32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_all_one_w_range35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_all_one_w_range37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_all_one_w_range39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_all_one_w_range41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_all_one_w_range43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_all_one_w_range45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_all_one_w_range47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_not_zero_w_range8w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_not_zero_w_range12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_not_zero_w_range15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_not_zero_w_range18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_not_zero_w_range21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_not_zero_w_range24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_not_zero_w_range27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_all_one_w_range559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_all_one_w_range565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_all_one_w_range570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_all_one_w_range575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_all_one_w_range580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_all_one_w_range585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_all_one_w_range590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_not_zero_w_range561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_not_zero_w_range567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_not_zero_w_range572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_not_zero_w_range577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_not_zero_w_range582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_not_zero_w_range587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_out_not_zero_w_range592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_result_w_range563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_result_w_range568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_result_w_range573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_result_w_range578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_result_w_range583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_result_w_range588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_result_w_range593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_value_wo_range129w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_w_exp_value_wo_range132w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_exp_value_wo_range131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range80w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range83w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_data_not_zero_w_range77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_prod_result_range424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_prod_result_range421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_prod_result_range418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_prod_result_range415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_prod_wo_range402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_all_ones_range491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_round_wi_range489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bits_range413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bits_range417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bits_range420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bits_range423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_xf_pre_2_wo_range183w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_w_xf_pre_wo_range177w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_clshift
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_SHIFTTYPE	:	STRING := "LOGICAL";
		LPM_WIDTH	:	NATURAL;
		LPM_WIDTHDIST	:	NATURAL;
		lpm_type	:	STRING := "lpm_clshift"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		direction	:	IN STD_LOGIC := '0';
		distance	:	IN STD_LOGIC_VECTOR(LPM_WIDTHDIST-1 DOWNTO 0);
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		underflow	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	loop0 : FOR i IN 0 TO 61 GENERATE 
		wire_w_lg_man_prod_shifted408w(i) <= man_prod_shifted(i) AND wire_w_man_prod_wo_range402w(0);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 61 GENERATE 
		wire_w_lg_man_prod_wire407w(i) <= man_prod_wire(i) AND wire_w_lg_w_man_prod_wo_range402w406w(0);
	END GENERATE loop1;
	wire_w_lg_underflow_w554w(0) <= underflow_w AND wire_w_lg_barrel_shifter_underflow553w(0);
	wire_w_lg_w_data_range10w34w(0) <= wire_w_data_range10w(0) AND wire_w_exp_data_all_one_w_range32w(0);
	wire_w_lg_w_data_range13w36w(0) <= wire_w_data_range13w(0) AND wire_w_exp_data_all_one_w_range35w(0);
	wire_w_lg_w_data_range16w38w(0) <= wire_w_data_range16w(0) AND wire_w_exp_data_all_one_w_range37w(0);
	wire_w_lg_w_data_range19w40w(0) <= wire_w_data_range19w(0) AND wire_w_exp_data_all_one_w_range39w(0);
	wire_w_lg_w_data_range22w42w(0) <= wire_w_data_range22w(0) AND wire_w_exp_data_all_one_w_range41w(0);
	wire_w_lg_w_data_range25w44w(0) <= wire_w_data_range25w(0) AND wire_w_exp_data_all_one_w_range43w(0);
	wire_w_lg_w_data_range28w46w(0) <= wire_w_data_range28w(0) AND wire_w_exp_data_all_one_w_range45w(0);
	wire_w_lg_w_exp_data_all_one_w_range47w119w(0) <= wire_w_exp_data_all_one_w_range47w(0) AND wire_w_lg_w_man_data_not_zero_w_range116w118w(0);
	wire_w_lg_w_exp_result_w_range563w564w(0) <= wire_w_exp_result_w_range563w(0) AND wire_w_exp_out_all_one_w_range559w(0);
	wire_w_lg_w_exp_result_w_range568w569w(0) <= wire_w_exp_result_w_range568w(0) AND wire_w_exp_out_all_one_w_range565w(0);
	wire_w_lg_w_exp_result_w_range573w574w(0) <= wire_w_exp_result_w_range573w(0) AND wire_w_exp_out_all_one_w_range570w(0);
	wire_w_lg_w_exp_result_w_range578w579w(0) <= wire_w_exp_result_w_range578w(0) AND wire_w_exp_out_all_one_w_range575w(0);
	wire_w_lg_w_exp_result_w_range583w584w(0) <= wire_w_exp_result_w_range583w(0) AND wire_w_exp_out_all_one_w_range580w(0);
	wire_w_lg_w_exp_result_w_range588w589w(0) <= wire_w_exp_result_w_range588w(0) AND wire_w_exp_out_all_one_w_range585w(0);
	wire_w_lg_w_exp_result_w_range593w594w(0) <= wire_w_exp_result_w_range593w(0) AND wire_w_exp_out_all_one_w_range590w(0);
	wire_w_lg_w_man_round_wi_range492w493w(0) <= wire_w_man_round_wi_range492w(0) AND wire_w_man_result_all_ones_range491w(0);
	wire_w_lg_w_man_round_wi_range495w496w(0) <= wire_w_man_round_wi_range495w(0) AND wire_w_man_result_all_ones_range494w(0);
	wire_w_lg_w_man_round_wi_range498w499w(0) <= wire_w_man_round_wi_range498w(0) AND wire_w_man_result_all_ones_range497w(0);
	wire_w_lg_w_man_round_wi_range501w502w(0) <= wire_w_man_round_wi_range501w(0) AND wire_w_man_result_all_ones_range500w(0);
	wire_w_lg_w_man_round_wi_range504w505w(0) <= wire_w_man_round_wi_range504w(0) AND wire_w_man_result_all_ones_range503w(0);
	wire_w_lg_w_man_round_wi_range507w508w(0) <= wire_w_man_round_wi_range507w(0) AND wire_w_man_result_all_ones_range506w(0);
	wire_w_lg_w_man_round_wi_range510w511w(0) <= wire_w_man_round_wi_range510w(0) AND wire_w_man_result_all_ones_range509w(0);
	wire_w_lg_w_man_round_wi_range513w514w(0) <= wire_w_man_round_wi_range513w(0) AND wire_w_man_result_all_ones_range512w(0);
	wire_w_lg_w_man_round_wi_range516w517w(0) <= wire_w_man_round_wi_range516w(0) AND wire_w_man_result_all_ones_range515w(0);
	wire_w_lg_w_man_round_wi_range519w520w(0) <= wire_w_man_round_wi_range519w(0) AND wire_w_man_result_all_ones_range518w(0);
	wire_w_lg_w_man_round_wi_range465w466w(0) <= wire_w_man_round_wi_range465w(0) AND wire_w_man_result_all_ones_range463w(0);
	wire_w_lg_w_man_round_wi_range522w523w(0) <= wire_w_man_round_wi_range522w(0) AND wire_w_man_result_all_ones_range521w(0);
	wire_w_lg_w_man_round_wi_range525w526w(0) <= wire_w_man_round_wi_range525w(0) AND wire_w_man_result_all_ones_range524w(0);
	wire_w_lg_w_man_round_wi_range528w529w(0) <= wire_w_man_round_wi_range528w(0) AND wire_w_man_result_all_ones_range527w(0);
	wire_w_lg_w_man_round_wi_range468w469w(0) <= wire_w_man_round_wi_range468w(0) AND wire_w_man_result_all_ones_range467w(0);
	wire_w_lg_w_man_round_wi_range471w472w(0) <= wire_w_man_round_wi_range471w(0) AND wire_w_man_result_all_ones_range470w(0);
	wire_w_lg_w_man_round_wi_range474w475w(0) <= wire_w_man_round_wi_range474w(0) AND wire_w_man_result_all_ones_range473w(0);
	wire_w_lg_w_man_round_wi_range477w478w(0) <= wire_w_man_round_wi_range477w(0) AND wire_w_man_result_all_ones_range476w(0);
	wire_w_lg_w_man_round_wi_range480w481w(0) <= wire_w_man_round_wi_range480w(0) AND wire_w_man_result_all_ones_range479w(0);
	wire_w_lg_w_man_round_wi_range483w484w(0) <= wire_w_man_round_wi_range483w(0) AND wire_w_man_result_all_ones_range482w(0);
	wire_w_lg_w_man_round_wi_range486w487w(0) <= wire_w_man_round_wi_range486w(0) AND wire_w_man_result_all_ones_range485w(0);
	wire_w_lg_w_man_round_wi_range489w490w(0) <= wire_w_man_round_wi_range489w(0) AND wire_w_man_result_all_ones_range488w(0);
	wire_w_lg_w_lg_w_lg_underflow_w554w555w556w(0) <= NOT wire_w_lg_w_lg_underflow_w554w555w(0);
	wire_w_lg_barrel_shifter_underflow553w(0) <= NOT barrel_shifter_underflow;
	wire_w_lg_input_is_infinity_wo443w(0) <= NOT input_is_infinity_wo;
	wire_w_lg_input_is_nan_wo442w(0) <= NOT input_is_nan_wo;
	wire_w_lg_input_is_zero_wo444w(0) <= NOT input_is_zero_wo;
	wire_w_lg_underflow_w454w(0) <= NOT underflow_w;
	wire_w_lg_w_man_data_not_zero_w_range116w118w(0) <= NOT wire_w_man_data_not_zero_w_range116w(0);
	wire_w_lg_w_man_prod_wo_range402w406w(0) <= NOT wire_w_man_prod_wo_range402w(0);
	wire_w_lg_w_lg_underflow_w554w555w(0) <= wire_w_lg_underflow_w554w(0) OR negative_infinity;
	wire_w_lg_w551w552w(0) <= wire_w551w(0) OR positive_infinity;
	wire_w_lg_w_lg_w_lg_w_lg_overflow_w536w537w538w539w(0) <= wire_w_lg_w_lg_w_lg_overflow_w536w537w538w(0) OR input_is_infinity_wo;
	wire_w551w(0) <= wire_w_lg_w_lg_barrel_shifter_underflow549w550w(0) OR nan_w;
	wire_w_lg_w_lg_w_lg_overflow_w536w537w538w(0) <= wire_w_lg_w_lg_overflow_w536w537w(0) OR input_is_zero_wo;
	wire_w_lg_w_lg_barrel_shifter_underflow549w550w(0) <= wire_w_lg_barrel_shifter_underflow549w(0) OR input_is_zero_wo;
	wire_w_lg_w_lg_overflow_w542w543w(0) <= wire_w_lg_overflow_w542w(0) OR positive_infinity;
	wire_w_lg_w_lg_overflow_w536w537w(0) <= wire_w_lg_overflow_w536w(0) OR nan_w;
	wire_w_lg_barrel_shifter_underflow549w(0) <= barrel_shifter_underflow OR overflow_w;
	wire_w_lg_distance_overflow447w(0) <= distance_overflow OR wire_exp_value_add_bias_w_lg_w_result_range445w446w(0);
	wire_w_lg_distance_overflow456w(0) <= distance_overflow OR wire_exp_value_add_bias_w_result_range445w(0);
	wire_w_lg_overflow_w542w(0) <= overflow_w OR nan_w;
	wire_w_lg_overflow_w536w(0) <= overflow_w OR underflow_w;
	wire_w_lg_w_data_range78w79w(0) <= wire_w_data_range78w(0) OR wire_w_man_data_not_zero_w_range77w(0);
	wire_w_lg_w_data_range81w82w(0) <= wire_w_data_range81w(0) OR wire_w_man_data_not_zero_w_range80w(0);
	wire_w_lg_w_data_range84w85w(0) <= wire_w_data_range84w(0) OR wire_w_man_data_not_zero_w_range83w(0);
	wire_w_lg_w_data_range87w88w(0) <= wire_w_data_range87w(0) OR wire_w_man_data_not_zero_w_range86w(0);
	wire_w_lg_w_data_range90w91w(0) <= wire_w_data_range90w(0) OR wire_w_man_data_not_zero_w_range89w(0);
	wire_w_lg_w_data_range93w94w(0) <= wire_w_data_range93w(0) OR wire_w_man_data_not_zero_w_range92w(0);
	wire_w_lg_w_data_range96w97w(0) <= wire_w_data_range96w(0) OR wire_w_man_data_not_zero_w_range95w(0);
	wire_w_lg_w_data_range99w100w(0) <= wire_w_data_range99w(0) OR wire_w_man_data_not_zero_w_range98w(0);
	wire_w_lg_w_data_range102w103w(0) <= wire_w_data_range102w(0) OR wire_w_man_data_not_zero_w_range101w(0);
	wire_w_lg_w_data_range105w106w(0) <= wire_w_data_range105w(0) OR wire_w_man_data_not_zero_w_range104w(0);
	wire_w_lg_w_data_range51w52w(0) <= wire_w_data_range51w(0) OR wire_w_man_data_not_zero_w_range49w(0);
	wire_w_lg_w_data_range108w109w(0) <= wire_w_data_range108w(0) OR wire_w_man_data_not_zero_w_range107w(0);
	wire_w_lg_w_data_range111w112w(0) <= wire_w_data_range111w(0) OR wire_w_man_data_not_zero_w_range110w(0);
	wire_w_lg_w_data_range114w115w(0) <= wire_w_data_range114w(0) OR wire_w_man_data_not_zero_w_range113w(0);
	wire_w_lg_w_data_range10w11w(0) <= wire_w_data_range10w(0) OR wire_w_exp_data_not_zero_w_range8w(0);
	wire_w_lg_w_data_range13w14w(0) <= wire_w_data_range13w(0) OR wire_w_exp_data_not_zero_w_range12w(0);
	wire_w_lg_w_data_range16w17w(0) <= wire_w_data_range16w(0) OR wire_w_exp_data_not_zero_w_range15w(0);
	wire_w_lg_w_data_range19w20w(0) <= wire_w_data_range19w(0) OR wire_w_exp_data_not_zero_w_range18w(0);
	wire_w_lg_w_data_range22w23w(0) <= wire_w_data_range22w(0) OR wire_w_exp_data_not_zero_w_range21w(0);
	wire_w_lg_w_data_range25w26w(0) <= wire_w_data_range25w(0) OR wire_w_exp_data_not_zero_w_range24w(0);
	wire_w_lg_w_data_range54w55w(0) <= wire_w_data_range54w(0) OR wire_w_man_data_not_zero_w_range53w(0);
	wire_w_lg_w_data_range28w29w(0) <= wire_w_data_range28w(0) OR wire_w_exp_data_not_zero_w_range27w(0);
	wire_w_lg_w_data_range57w58w(0) <= wire_w_data_range57w(0) OR wire_w_man_data_not_zero_w_range56w(0);
	wire_w_lg_w_data_range60w61w(0) <= wire_w_data_range60w(0) OR wire_w_man_data_not_zero_w_range59w(0);
	wire_w_lg_w_data_range63w64w(0) <= wire_w_data_range63w(0) OR wire_w_man_data_not_zero_w_range62w(0);
	wire_w_lg_w_data_range66w67w(0) <= wire_w_data_range66w(0) OR wire_w_man_data_not_zero_w_range65w(0);
	wire_w_lg_w_data_range69w70w(0) <= wire_w_data_range69w(0) OR wire_w_man_data_not_zero_w_range68w(0);
	wire_w_lg_w_data_range72w73w(0) <= wire_w_data_range72w(0) OR wire_w_man_data_not_zero_w_range71w(0);
	wire_w_lg_w_data_range75w76w(0) <= wire_w_data_range75w(0) OR wire_w_man_data_not_zero_w_range74w(0);
	wire_w_lg_w_exp_result_w_range563w566w(0) <= wire_w_exp_result_w_range563w(0) OR wire_w_exp_out_not_zero_w_range561w(0);
	wire_w_lg_w_exp_result_w_range568w571w(0) <= wire_w_exp_result_w_range568w(0) OR wire_w_exp_out_not_zero_w_range567w(0);
	wire_w_lg_w_exp_result_w_range573w576w(0) <= wire_w_exp_result_w_range573w(0) OR wire_w_exp_out_not_zero_w_range572w(0);
	wire_w_lg_w_exp_result_w_range578w581w(0) <= wire_w_exp_result_w_range578w(0) OR wire_w_exp_out_not_zero_w_range577w(0);
	wire_w_lg_w_exp_result_w_range583w586w(0) <= wire_w_exp_result_w_range583w(0) OR wire_w_exp_out_not_zero_w_range582w(0);
	wire_w_lg_w_exp_result_w_range588w591w(0) <= wire_w_exp_result_w_range588w(0) OR wire_w_exp_out_not_zero_w_range587w(0);
	wire_w_lg_w_exp_result_w_range593w595w(0) <= wire_w_exp_result_w_range593w(0) OR wire_w_exp_out_not_zero_w_range592w(0);
	wire_w_lg_w_man_prod_result_range424w425w(0) <= wire_w_man_prod_result_range424w(0) OR wire_w_sticky_bits_range423w(0);
	wire_w_lg_w_man_prod_result_range421w422w(0) <= wire_w_man_prod_result_range421w(0) OR wire_w_sticky_bits_range420w(0);
	wire_w_lg_w_man_prod_result_range418w419w(0) <= wire_w_man_prod_result_range418w(0) OR wire_w_sticky_bits_range417w(0);
	wire_w_lg_w_man_prod_result_range415w416w(0) <= wire_w_man_prod_result_range415w(0) OR wire_w_sticky_bits_range413w(0);
	aclr <= '0';
	addr_val_more_than_one <= "10111";
	barrel_shifter_data <= ( "00000000" & "1" & fraction_wo & "000000");
	barrel_shifter_distance <= wire_exp_value_selecta_dataout;
	barrel_shifter_underflow <= barrel_shifter_underflow_dffe2_15_pipes14;
	barrel_shifter_underflow_wi <= (wire_underflow_compare_agb AND exp_value_wo(8));
	clk_en <= '1';
	distance_overflow <= distance_overflow_dffe2_15_pipes14;
	distance_overflow_val_w <= "00000110";
	distance_overflow_wi <= (wire_distance_overflow_comp_agb AND (NOT exp_value_wo(8)));
	exp_bias <= "01111111";
	exp_bias_all_ones_w <= (OTHERS => '1');
	exp_data_all_one_w <= ( wire_w_lg_w_data_range28w46w & wire_w_lg_w_data_range25w44w & wire_w_lg_w_data_range22w42w & wire_w_lg_w_data_range19w40w & wire_w_lg_w_data_range16w38w & wire_w_lg_w_data_range13w36w & wire_w_lg_w_data_range10w34w & data(23));
	exp_data_not_zero_w <= ( wire_w_lg_w_data_range28w29w & wire_w_lg_w_data_range25w26w & wire_w_lg_w_data_range22w23w & wire_w_lg_w_data_range19w20w & wire_w_lg_w_data_range16w17w & wire_w_lg_w_data_range13w14w & wire_w_lg_w_data_range10w11w & data(23));
	exp_invert <= (xi_exp_value XOR exp_bias_all_ones_w);
	exp_one <= ( wire_w_lg_w_lg_overflow_w542w543w & "1111111");
	exp_out_all_one_w <= ( wire_w_lg_w_exp_result_w_range593w594w & wire_w_lg_w_exp_result_w_range588w589w & wire_w_lg_w_exp_result_w_range583w584w & wire_w_lg_w_exp_result_w_range578w579w & wire_w_lg_w_exp_result_w_range573w574w & wire_w_lg_w_exp_result_w_range568w569w & wire_w_lg_w_exp_result_w_range563w564w & exp_result_w(0));
	exp_out_not_zero_w <= ( wire_w_lg_w_exp_result_w_range593w595w & wire_w_lg_w_exp_result_w_range588w591w & wire_w_lg_w_exp_result_w_range583w586w & wire_w_lg_w_exp_result_w_range578w581w & wire_w_lg_w_exp_result_w_range573w576w & wire_w_lg_w_exp_result_w_range568w571w & wire_w_lg_w_exp_result_w_range563w566w & exp_result_w(0));
	exp_result_out <= wire_exp_result_mux_prea_w_lg_dataout557w;
	exp_result_w <= wire_exp_value_man_over_result(7 DOWNTO 0);
	exp_value <= wire_exp_minus_bias_result;
	exp_value_wi <= exp_value;
	exp_value_wo <= exp_value_dffe1;
	exp_w <= data(30 DOWNTO 23);
	extra_ln2 <= ((NOT xf_pre(37)) AND sign_dffe8);
	fraction <= ( data(22 DOWNTO 0));
	fraction_wi <= fraction;
	fraction_wo <= fraction_dffe1;
	gnd_w <= '0';
	guard_bit <= man_prod_result(35);
	input_is_infinity_wi <= wire_w_lg_w_exp_data_all_one_w_range47w119w(0);
	input_is_infinity_wo <= input_is_infinity_16_pipes15;
	input_is_nan_wi <= (exp_data_all_one_w(7) AND man_data_not_zero_w(22));
	input_is_nan_wo <= input_is_nan_16_pipes15;
	input_is_zero_wi <= (NOT exp_data_not_zero_w(7));
	input_is_zero_wo <= input_is_zero_16_pipes15;
	ln2_w <= "10110001011100100001011111110111110100";
	man_data_not_zero_w <= ( wire_w_lg_w_data_range114w115w & wire_w_lg_w_data_range111w112w & wire_w_lg_w_data_range108w109w & wire_w_lg_w_data_range105w106w & wire_w_lg_w_data_range102w103w & wire_w_lg_w_data_range99w100w & wire_w_lg_w_data_range96w97w & wire_w_lg_w_data_range93w94w & wire_w_lg_w_data_range90w91w & wire_w_lg_w_data_range87w88w & wire_w_lg_w_data_range84w85w & wire_w_lg_w_data_range81w82w & wire_w_lg_w_data_range78w79w & wire_w_lg_w_data_range75w76w & wire_w_lg_w_data_range72w73w & wire_w_lg_w_data_range69w70w & wire_w_lg_w_data_range66w67w & wire_w_lg_w_data_range63w64w & wire_w_lg_w_data_range60w61w & wire_w_lg_w_data_range57w58w & wire_w_lg_w_data_range54w55w & wire_w_lg_w_data_range51w52w & data(0));
	man_overflow <= (round_up AND man_result_all_ones(22));
	man_overflow_wi <= man_overflow;
	man_overflow_wo <= man_overflow_dffe15;
	man_prod_result <= (wire_w_lg_man_prod_shifted408w OR wire_w_lg_man_prod_wire407w);
	man_prod_shifted <= ( gnd_w & man_prod_wo(61 DOWNTO 1));
	man_prod_wi <= wire_man_prod_result;
	man_prod_wire <= man_prod_wo;
	man_prod_wo <= man_prod_dffe14;
	man_result_all_ones <= ( wire_w_lg_w_man_round_wi_range528w529w & wire_w_lg_w_man_round_wi_range525w526w & wire_w_lg_w_man_round_wi_range522w523w & wire_w_lg_w_man_round_wi_range519w520w & wire_w_lg_w_man_round_wi_range516w517w & wire_w_lg_w_man_round_wi_range513w514w & wire_w_lg_w_man_round_wi_range510w511w & wire_w_lg_w_man_round_wi_range507w508w & wire_w_lg_w_man_round_wi_range504w505w & wire_w_lg_w_man_round_wi_range501w502w & wire_w_lg_w_man_round_wi_range498w499w & wire_w_lg_w_man_round_wi_range495w496w & wire_w_lg_w_man_round_wi_range492w493w & wire_w_lg_w_man_round_wi_range489w490w & wire_w_lg_w_man_round_wi_range486w487w & wire_w_lg_w_man_round_wi_range483w484w & wire_w_lg_w_man_round_wi_range480w481w & wire_w_lg_w_man_round_wi_range477w478w & wire_w_lg_w_man_round_wi_range474w475w & wire_w_lg_w_man_round_wi_range471w472w & wire_w_lg_w_man_round_wi_range468w469w & wire_w_lg_w_man_round_wi_range465w466w & man_round_wi(0));
	man_result_w <= wire_man_result_muxa_dataout;
	man_round_wi <= man_prod_result(57 DOWNTO 35);
	man_round_wo <= man_round_dffe15;
	nan_w <= input_is_nan_wo;
	negative_infinity <= (sign_dffe15 AND input_is_infinity_wo);
	one_over_ln2_w <= "101110001";
	overflow_w <= (((wire_sign_dffe_w_lg_q434w(0) AND ((wire_w_lg_distance_overflow456w(0) OR exp_out_all_one_w(7)) OR wire_exp_value_man_over_result(8))) AND wire_w_lg_underflow_w454w(0)) AND wire_w_lg_input_is_nan_wo442w(0));
	positive_infinity <= (wire_sign_dffe_w_lg_q434w(0) AND input_is_infinity_wo);
	result <= ( "0" & result_pipe_wo);
	result_pipe_wi <= ( exp_result_out & man_result_w);
	result_pipe_wo <= result_pipe_dffe16;
	result_underflow_w <= ((NOT exp_out_not_zero_w(7)) AND wire_exp_value_man_over_w_lg_w_lg_w_lg_w_result_range435w436w437w438w(0));
	round_bit <= man_prod_result(34);
	round_up <= (round_bit AND (guard_bit OR sticky_bits(4)));
	round_up_wi <= round_up;
	round_up_wo <= round_up_dffe15;
	shifted_value <= (tbl1_compare_wo OR man_prod_wo(59));
	sign_w <= data(31);
	sticky_bits <= ( wire_w_lg_w_man_prod_result_range424w425w & wire_w_lg_w_man_prod_result_range421w422w & wire_w_lg_w_man_prod_result_range418w419w & wire_w_lg_w_man_prod_result_range415w416w & man_prod_result(33));
	table_one_data <= ( "10101000100111100001011100110110" & "10100011011011100000001001111010" & "10011110011001101100101000011001" & "10011001100001110010110000111101" & "10010100110011011111000011111001" & "10010000001110011110100111111000" & "10001011110010011111001000110010" & "10000111011111001110110110100011" & "10000011010100011100100100000011" & "11111110100011101111001100001100" & "11110110101110011111100100100000" & "11101111001000101010111011111100" & "11100111110001110010111011000010" & "11100000101001011010000110001001" & "11011001101111000011111011100100" & "11010011000010010100110001110000" & "11001100100010110001110101101010" & "11000110010000000001001000111011" & "11000000001001101001100000011010" & "10111010001111010010100010011110" & "10110100100000100100100101100101" & "10101110111101001000101110110000" & "10101001100100101000110000000110" & "10100100010110101111000111100001" & "10011111010011000110111101010101" & "10011010011001011100000010111000" & "10010101101001011010110001011001" & "10010001000010110000001000101101" & "10001100100101001001101110000011" & "10001000010000010101101010111011" & "10000100000100000010101100000000" & "10000000000000000000000000000000");
	table_one_out <= wire_table_one_result;
	table_three_data <= ( "111110000001111000001" & "111100000001110000100" & "111010000001101001001" & "111000000001100010000" & "110110000001011011001" & "110100000001010100100" & "110010000001001110001" & "110000000001001000000" & "101110000001000010001" & "101100000000111100100" & "101010000000110111001" & "101000000000110010000" & "100110000000101101001" & "100100000000101000100" & "100010000000100100001" & "100000000000100000000" & "011110000000011100001" & "011100000000011000100" & "011010000000010101001" & "011000000000010010000" & "010110000000001111001" & "010100000000001100100" & "010010000000001010001" & "010000000000001000000" & "001110000000000110001" & "001100000000000100100" & "001010000000000011001" & "001000000000000010000" & "000110000000000001001" & "000100000000000000100" & "000010000000000000001" & "000000000000000000000");
	table_three_out <= ( "1" & "0000000000" & table_three_out_tmp);
	table_three_out_tmp <= wire_table_three_result;
	table_two_data <= ( "11111011110010101100010101" & "11110011100011001101101010" & "11101011010100001111111011" & "11100011000101110011000111" & "11011010110111110111001100" & "11010010101010011100001000" & "11001010011101100001111000" & "11000010010001001000011011" & "10111010000101001111101110" & "10110001111001110111110000" & "10101001101111000000011110" & "10100001100100101001110111" & "10011001011010110011111000" & "10010001010001011110100000" & "10001001001000101001101100" & "10000001000000010101011010" & "01111000111000100001101001" & "01110000110001001110010101" & "01101000101010011011011110" & "01100000100100001001000001" & "01011000011110010110111100" & "01010000011001000101001110" & "01001000010100010011110011" & "01000000010000000010101011" & "00111000001100010001110010" & "00110000001001000001001000" & "00101000000110010000101001" & "00100000000100000000010101" & "00011000000010010000001001" & "00010000000001000000000010" & "00001000000000010000000000" & "00000000000000000000000000");
	table_two_out <= ( "1" & "00000" & table_two_out_tmp);
	table_two_out_tmp <= wire_table_two_result;
	tbl1_compare_wi <= wire_tbl1_compare_ageb;
	tbl1_compare_wo <= tbl1_compare_dffe11_4_pipes3;
	tbl1_tbl2_prod_wi <= wire_tbl1_tbl2_prod_result(63 DOWNTO 33);
	tbl1_tbl2_prod_wo <= tbl1_tbl2_prod_dffe12;
	tbl3_taylor_prod_wi <= wire_tbl3_taylor_prod_result(61 DOWNTO 31);
	tbl3_taylor_prod_wo <= tbl3_taylor_prod_dffe12;
	underflow_compare_val_w <= "00011101";
	underflow_w <= (((((result_underflow_w OR barrel_shifter_underflow) OR wire_sign_dffe_w_lg_q448w(0)) AND wire_w_lg_input_is_zero_wo444w(0)) AND wire_w_lg_input_is_infinity_wo443w(0)) AND wire_w_lg_input_is_nan_wo442w(0));
	x_fixed <= wire_rbarrel_shift_result;
	xf <= wire_xf_muxa_dataout;
	xf_pre <= wire_x_fixed_minus_xiln2_result;
	xf_pre_2_wi <= xf_pre_wo;
	xf_pre_2_wo <= xf_pre_2_dffe10;
	xf_pre_wi <= xf_pre;
	xf_pre_wo <= xf_pre_dffe9;
	xi_exp_value <= xi_prod_wo(18 DOWNTO 11);
	xi_exp_value_wi <= xi_exp_value;
	xi_exp_value_wo <= xi_exp_value_dffe4;
	xi_ln2_prod_wi <= wire_xi_ln2_prod_result;
	xi_ln2_prod_wo <= xi_ln2_prod_dffe7;
	xi_prod_wi <= wire_xi_prod_result;
	xi_prod_wo <= xi_prod_dffe3;
	wire_w_data_range78w(0) <= data(10);
	wire_w_data_range81w(0) <= data(11);
	wire_w_data_range84w(0) <= data(12);
	wire_w_data_range87w(0) <= data(13);
	wire_w_data_range90w(0) <= data(14);
	wire_w_data_range93w(0) <= data(15);
	wire_w_data_range96w(0) <= data(16);
	wire_w_data_range99w(0) <= data(17);
	wire_w_data_range102w(0) <= data(18);
	wire_w_data_range105w(0) <= data(19);
	wire_w_data_range51w(0) <= data(1);
	wire_w_data_range108w(0) <= data(20);
	wire_w_data_range111w(0) <= data(21);
	wire_w_data_range114w(0) <= data(22);
	wire_w_data_range10w(0) <= data(24);
	wire_w_data_range13w(0) <= data(25);
	wire_w_data_range16w(0) <= data(26);
	wire_w_data_range19w(0) <= data(27);
	wire_w_data_range22w(0) <= data(28);
	wire_w_data_range25w(0) <= data(29);
	wire_w_data_range54w(0) <= data(2);
	wire_w_data_range28w(0) <= data(30);
	wire_w_data_range57w(0) <= data(3);
	wire_w_data_range60w(0) <= data(4);
	wire_w_data_range63w(0) <= data(5);
	wire_w_data_range66w(0) <= data(6);
	wire_w_data_range69w(0) <= data(7);
	wire_w_data_range72w(0) <= data(8);
	wire_w_data_range75w(0) <= data(9);
	wire_w_exp_data_all_one_w_range32w(0) <= exp_data_all_one_w(0);
	wire_w_exp_data_all_one_w_range35w(0) <= exp_data_all_one_w(1);
	wire_w_exp_data_all_one_w_range37w(0) <= exp_data_all_one_w(2);
	wire_w_exp_data_all_one_w_range39w(0) <= exp_data_all_one_w(3);
	wire_w_exp_data_all_one_w_range41w(0) <= exp_data_all_one_w(4);
	wire_w_exp_data_all_one_w_range43w(0) <= exp_data_all_one_w(5);
	wire_w_exp_data_all_one_w_range45w(0) <= exp_data_all_one_w(6);
	wire_w_exp_data_all_one_w_range47w(0) <= exp_data_all_one_w(7);
	wire_w_exp_data_not_zero_w_range8w(0) <= exp_data_not_zero_w(0);
	wire_w_exp_data_not_zero_w_range12w(0) <= exp_data_not_zero_w(1);
	wire_w_exp_data_not_zero_w_range15w(0) <= exp_data_not_zero_w(2);
	wire_w_exp_data_not_zero_w_range18w(0) <= exp_data_not_zero_w(3);
	wire_w_exp_data_not_zero_w_range21w(0) <= exp_data_not_zero_w(4);
	wire_w_exp_data_not_zero_w_range24w(0) <= exp_data_not_zero_w(5);
	wire_w_exp_data_not_zero_w_range27w(0) <= exp_data_not_zero_w(6);
	wire_w_exp_out_all_one_w_range559w(0) <= exp_out_all_one_w(0);
	wire_w_exp_out_all_one_w_range565w(0) <= exp_out_all_one_w(1);
	wire_w_exp_out_all_one_w_range570w(0) <= exp_out_all_one_w(2);
	wire_w_exp_out_all_one_w_range575w(0) <= exp_out_all_one_w(3);
	wire_w_exp_out_all_one_w_range580w(0) <= exp_out_all_one_w(4);
	wire_w_exp_out_all_one_w_range585w(0) <= exp_out_all_one_w(5);
	wire_w_exp_out_all_one_w_range590w(0) <= exp_out_all_one_w(6);
	wire_w_exp_out_not_zero_w_range561w(0) <= exp_out_not_zero_w(0);
	wire_w_exp_out_not_zero_w_range567w(0) <= exp_out_not_zero_w(1);
	wire_w_exp_out_not_zero_w_range572w(0) <= exp_out_not_zero_w(2);
	wire_w_exp_out_not_zero_w_range577w(0) <= exp_out_not_zero_w(3);
	wire_w_exp_out_not_zero_w_range582w(0) <= exp_out_not_zero_w(4);
	wire_w_exp_out_not_zero_w_range587w(0) <= exp_out_not_zero_w(5);
	wire_w_exp_out_not_zero_w_range592w(0) <= exp_out_not_zero_w(6);
	wire_w_exp_result_w_range563w(0) <= exp_result_w(1);
	wire_w_exp_result_w_range568w(0) <= exp_result_w(2);
	wire_w_exp_result_w_range573w(0) <= exp_result_w(3);
	wire_w_exp_result_w_range578w(0) <= exp_result_w(4);
	wire_w_exp_result_w_range583w(0) <= exp_result_w(5);
	wire_w_exp_result_w_range588w(0) <= exp_result_w(6);
	wire_w_exp_result_w_range593w(0) <= exp_result_w(7);
	wire_w_exp_value_wo_range129w <= exp_value_wo(5 DOWNTO 0);
	wire_w_exp_value_wo_range132w <= exp_value_wo(7 DOWNTO 0);
	wire_w_exp_value_wo_range131w(0) <= exp_value_wo(8);
	wire_w_man_data_not_zero_w_range49w(0) <= man_data_not_zero_w(0);
	wire_w_man_data_not_zero_w_range80w(0) <= man_data_not_zero_w(10);
	wire_w_man_data_not_zero_w_range83w(0) <= man_data_not_zero_w(11);
	wire_w_man_data_not_zero_w_range86w(0) <= man_data_not_zero_w(12);
	wire_w_man_data_not_zero_w_range89w(0) <= man_data_not_zero_w(13);
	wire_w_man_data_not_zero_w_range92w(0) <= man_data_not_zero_w(14);
	wire_w_man_data_not_zero_w_range95w(0) <= man_data_not_zero_w(15);
	wire_w_man_data_not_zero_w_range98w(0) <= man_data_not_zero_w(16);
	wire_w_man_data_not_zero_w_range101w(0) <= man_data_not_zero_w(17);
	wire_w_man_data_not_zero_w_range104w(0) <= man_data_not_zero_w(18);
	wire_w_man_data_not_zero_w_range107w(0) <= man_data_not_zero_w(19);
	wire_w_man_data_not_zero_w_range53w(0) <= man_data_not_zero_w(1);
	wire_w_man_data_not_zero_w_range110w(0) <= man_data_not_zero_w(20);
	wire_w_man_data_not_zero_w_range113w(0) <= man_data_not_zero_w(21);
	wire_w_man_data_not_zero_w_range116w(0) <= man_data_not_zero_w(22);
	wire_w_man_data_not_zero_w_range56w(0) <= man_data_not_zero_w(2);
	wire_w_man_data_not_zero_w_range59w(0) <= man_data_not_zero_w(3);
	wire_w_man_data_not_zero_w_range62w(0) <= man_data_not_zero_w(4);
	wire_w_man_data_not_zero_w_range65w(0) <= man_data_not_zero_w(5);
	wire_w_man_data_not_zero_w_range68w(0) <= man_data_not_zero_w(6);
	wire_w_man_data_not_zero_w_range71w(0) <= man_data_not_zero_w(7);
	wire_w_man_data_not_zero_w_range74w(0) <= man_data_not_zero_w(8);
	wire_w_man_data_not_zero_w_range77w(0) <= man_data_not_zero_w(9);
	wire_w_man_prod_result_range424w(0) <= man_prod_result(29);
	wire_w_man_prod_result_range421w(0) <= man_prod_result(30);
	wire_w_man_prod_result_range418w(0) <= man_prod_result(31);
	wire_w_man_prod_result_range415w(0) <= man_prod_result(32);
	wire_w_man_prod_wo_range402w(0) <= man_prod_wo(59);
	wire_w_man_result_all_ones_range463w(0) <= man_result_all_ones(0);
	wire_w_man_result_all_ones_range494w(0) <= man_result_all_ones(10);
	wire_w_man_result_all_ones_range497w(0) <= man_result_all_ones(11);
	wire_w_man_result_all_ones_range500w(0) <= man_result_all_ones(12);
	wire_w_man_result_all_ones_range503w(0) <= man_result_all_ones(13);
	wire_w_man_result_all_ones_range506w(0) <= man_result_all_ones(14);
	wire_w_man_result_all_ones_range509w(0) <= man_result_all_ones(15);
	wire_w_man_result_all_ones_range512w(0) <= man_result_all_ones(16);
	wire_w_man_result_all_ones_range515w(0) <= man_result_all_ones(17);
	wire_w_man_result_all_ones_range518w(0) <= man_result_all_ones(18);
	wire_w_man_result_all_ones_range521w(0) <= man_result_all_ones(19);
	wire_w_man_result_all_ones_range467w(0) <= man_result_all_ones(1);
	wire_w_man_result_all_ones_range524w(0) <= man_result_all_ones(20);
	wire_w_man_result_all_ones_range527w(0) <= man_result_all_ones(21);
	wire_w_man_result_all_ones_range470w(0) <= man_result_all_ones(2);
	wire_w_man_result_all_ones_range473w(0) <= man_result_all_ones(3);
	wire_w_man_result_all_ones_range476w(0) <= man_result_all_ones(4);
	wire_w_man_result_all_ones_range479w(0) <= man_result_all_ones(5);
	wire_w_man_result_all_ones_range482w(0) <= man_result_all_ones(6);
	wire_w_man_result_all_ones_range485w(0) <= man_result_all_ones(7);
	wire_w_man_result_all_ones_range488w(0) <= man_result_all_ones(8);
	wire_w_man_result_all_ones_range491w(0) <= man_result_all_ones(9);
	wire_w_man_round_wi_range492w(0) <= man_round_wi(10);
	wire_w_man_round_wi_range495w(0) <= man_round_wi(11);
	wire_w_man_round_wi_range498w(0) <= man_round_wi(12);
	wire_w_man_round_wi_range501w(0) <= man_round_wi(13);
	wire_w_man_round_wi_range504w(0) <= man_round_wi(14);
	wire_w_man_round_wi_range507w(0) <= man_round_wi(15);
	wire_w_man_round_wi_range510w(0) <= man_round_wi(16);
	wire_w_man_round_wi_range513w(0) <= man_round_wi(17);
	wire_w_man_round_wi_range516w(0) <= man_round_wi(18);
	wire_w_man_round_wi_range519w(0) <= man_round_wi(19);
	wire_w_man_round_wi_range465w(0) <= man_round_wi(1);
	wire_w_man_round_wi_range522w(0) <= man_round_wi(20);
	wire_w_man_round_wi_range525w(0) <= man_round_wi(21);
	wire_w_man_round_wi_range528w(0) <= man_round_wi(22);
	wire_w_man_round_wi_range468w(0) <= man_round_wi(2);
	wire_w_man_round_wi_range471w(0) <= man_round_wi(3);
	wire_w_man_round_wi_range474w(0) <= man_round_wi(4);
	wire_w_man_round_wi_range477w(0) <= man_round_wi(5);
	wire_w_man_round_wi_range480w(0) <= man_round_wi(6);
	wire_w_man_round_wi_range483w(0) <= man_round_wi(7);
	wire_w_man_round_wi_range486w(0) <= man_round_wi(8);
	wire_w_man_round_wi_range489w(0) <= man_round_wi(9);
	wire_w_sticky_bits_range413w(0) <= sticky_bits(0);
	wire_w_sticky_bits_range417w(0) <= sticky_bits(1);
	wire_w_sticky_bits_range420w(0) <= sticky_bits(2);
	wire_w_sticky_bits_range423w(0) <= sticky_bits(3);
	wire_w_xf_pre_2_wo_range183w <= xf_pre_2_wo(30 DOWNTO 0);
	wire_w_xf_pre_wo_range177w <= xf_pre_wo(30 DOWNTO 0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_15_pipes0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_15_pipes0 <= barrel_shifter_underflow_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_15_pipes1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_15_pipes1 <= barrel_shifter_underflow_dffe2_15_pipes0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_15_pipes2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_15_pipes2 <= barrel_shifter_underflow_dffe2_15_pipes1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_15_pipes3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_15_pipes3 <= barrel_shifter_underflow_dffe2_15_pipes2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_15_pipes4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_15_pipes4 <= barrel_shifter_underflow_dffe2_15_pipes3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_15_pipes5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_15_pipes5 <= barrel_shifter_underflow_dffe2_15_pipes4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_15_pipes6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_15_pipes6 <= barrel_shifter_underflow_dffe2_15_pipes5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_15_pipes7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_15_pipes7 <= barrel_shifter_underflow_dffe2_15_pipes6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_15_pipes8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_15_pipes8 <= barrel_shifter_underflow_dffe2_15_pipes7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_15_pipes9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_15_pipes9 <= barrel_shifter_underflow_dffe2_15_pipes8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_15_pipes10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_15_pipes10 <= barrel_shifter_underflow_dffe2_15_pipes9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_15_pipes11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_15_pipes11 <= barrel_shifter_underflow_dffe2_15_pipes10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_15_pipes12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_15_pipes12 <= barrel_shifter_underflow_dffe2_15_pipes11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_15_pipes13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_15_pipes13 <= barrel_shifter_underflow_dffe2_15_pipes12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN barrel_shifter_underflow_dffe2_15_pipes14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN barrel_shifter_underflow_dffe2_15_pipes14 <= barrel_shifter_underflow_dffe2_15_pipes13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_15_pipes0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_15_pipes0 <= distance_overflow_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_15_pipes1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_15_pipes1 <= distance_overflow_dffe2_15_pipes0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_15_pipes2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_15_pipes2 <= distance_overflow_dffe2_15_pipes1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_15_pipes3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_15_pipes3 <= distance_overflow_dffe2_15_pipes2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_15_pipes4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_15_pipes4 <= distance_overflow_dffe2_15_pipes3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_15_pipes5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_15_pipes5 <= distance_overflow_dffe2_15_pipes4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_15_pipes6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_15_pipes6 <= distance_overflow_dffe2_15_pipes5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_15_pipes7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_15_pipes7 <= distance_overflow_dffe2_15_pipes6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_15_pipes8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_15_pipes8 <= distance_overflow_dffe2_15_pipes7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_15_pipes9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_15_pipes9 <= distance_overflow_dffe2_15_pipes8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_15_pipes10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_15_pipes10 <= distance_overflow_dffe2_15_pipes9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_15_pipes11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_15_pipes11 <= distance_overflow_dffe2_15_pipes10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_15_pipes12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_15_pipes12 <= distance_overflow_dffe2_15_pipes11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_15_pipes13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_15_pipes13 <= distance_overflow_dffe2_15_pipes12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN distance_overflow_dffe2_15_pipes14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN distance_overflow_dffe2_15_pipes14 <= distance_overflow_dffe2_15_pipes13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_0 <= wire_exp_value_b4_biasa_dataout;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_1 <= exp_value_b4_bias_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_10 <= exp_value_b4_bias_dffe_9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_2 <= exp_value_b4_bias_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_3 <= exp_value_b4_bias_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_4 <= exp_value_b4_bias_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_5 <= exp_value_b4_bias_dffe_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_6 <= exp_value_b4_bias_dffe_5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_7 <= exp_value_b4_bias_dffe_6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_8 <= exp_value_b4_bias_dffe_7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_b4_bias_dffe_9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_b4_bias_dffe_9 <= exp_value_b4_bias_dffe_8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_value_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_value_dffe1 <= exp_value_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN extra_ln2_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN extra_ln2_dffe_0 <= extra_ln2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN extra_ln2_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN extra_ln2_dffe_1 <= extra_ln2_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN extra_ln2_dffe_2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN extra_ln2_dffe_2 <= extra_ln2_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN extra_ln2_dffe_3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN extra_ln2_dffe_3 <= extra_ln2_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN extra_ln2_dffe_4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN extra_ln2_dffe_4 <= extra_ln2_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN extra_ln2_dffe_5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN extra_ln2_dffe_5 <= extra_ln2_dffe_4;
			END IF;
		END IF;
	END PROCESS;
	wire_extra_ln2_dffe_5_w_lg_q157w(0) <= NOT extra_ln2_dffe_5;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN fraction_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN fraction_dffe1 <= fraction_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_16_pipes0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_16_pipes0 <= input_is_infinity_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_16_pipes1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_16_pipes1 <= input_is_infinity_16_pipes0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_16_pipes2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_16_pipes2 <= input_is_infinity_16_pipes1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_16_pipes3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_16_pipes3 <= input_is_infinity_16_pipes2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_16_pipes4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_16_pipes4 <= input_is_infinity_16_pipes3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_16_pipes5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_16_pipes5 <= input_is_infinity_16_pipes4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_16_pipes6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_16_pipes6 <= input_is_infinity_16_pipes5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_16_pipes7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_16_pipes7 <= input_is_infinity_16_pipes6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_16_pipes8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_16_pipes8 <= input_is_infinity_16_pipes7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_16_pipes9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_16_pipes9 <= input_is_infinity_16_pipes8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_16_pipes10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_16_pipes10 <= input_is_infinity_16_pipes9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_16_pipes11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_16_pipes11 <= input_is_infinity_16_pipes10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_16_pipes12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_16_pipes12 <= input_is_infinity_16_pipes11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_16_pipes13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_16_pipes13 <= input_is_infinity_16_pipes12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_16_pipes14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_16_pipes14 <= input_is_infinity_16_pipes13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_16_pipes15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_16_pipes15 <= input_is_infinity_16_pipes14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_16_pipes0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_16_pipes0 <= input_is_nan_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_16_pipes1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_16_pipes1 <= input_is_nan_16_pipes0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_16_pipes2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_16_pipes2 <= input_is_nan_16_pipes1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_16_pipes3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_16_pipes3 <= input_is_nan_16_pipes2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_16_pipes4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_16_pipes4 <= input_is_nan_16_pipes3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_16_pipes5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_16_pipes5 <= input_is_nan_16_pipes4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_16_pipes6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_16_pipes6 <= input_is_nan_16_pipes5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_16_pipes7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_16_pipes7 <= input_is_nan_16_pipes6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_16_pipes8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_16_pipes8 <= input_is_nan_16_pipes7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_16_pipes9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_16_pipes9 <= input_is_nan_16_pipes8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_16_pipes10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_16_pipes10 <= input_is_nan_16_pipes9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_16_pipes11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_16_pipes11 <= input_is_nan_16_pipes10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_16_pipes12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_16_pipes12 <= input_is_nan_16_pipes11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_16_pipes13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_16_pipes13 <= input_is_nan_16_pipes12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_16_pipes14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_16_pipes14 <= input_is_nan_16_pipes13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_16_pipes15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_16_pipes15 <= input_is_nan_16_pipes14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_16_pipes0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_16_pipes0 <= input_is_zero_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_16_pipes1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_16_pipes1 <= input_is_zero_16_pipes0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_16_pipes2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_16_pipes2 <= input_is_zero_16_pipes1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_16_pipes3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_16_pipes3 <= input_is_zero_16_pipes2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_16_pipes4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_16_pipes4 <= input_is_zero_16_pipes3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_16_pipes5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_16_pipes5 <= input_is_zero_16_pipes4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_16_pipes6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_16_pipes6 <= input_is_zero_16_pipes5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_16_pipes7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_16_pipes7 <= input_is_zero_16_pipes6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_16_pipes8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_16_pipes8 <= input_is_zero_16_pipes7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_16_pipes9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_16_pipes9 <= input_is_zero_16_pipes8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_16_pipes10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_16_pipes10 <= input_is_zero_16_pipes9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_16_pipes11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_16_pipes11 <= input_is_zero_16_pipes10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_16_pipes12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_16_pipes12 <= input_is_zero_16_pipes11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_16_pipes13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_16_pipes13 <= input_is_zero_16_pipes12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_16_pipes14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_16_pipes14 <= input_is_zero_16_pipes13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_16_pipes15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_16_pipes15 <= input_is_zero_16_pipes14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_overflow_dffe15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_overflow_dffe15 <= man_overflow_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_prod_dffe14 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_prod_dffe14 <= man_prod_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_round_dffe15 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_round_dffe15 <= man_round_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN result_pipe_dffe16 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN result_pipe_dffe16 <= result_pipe_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN round_up_dffe15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN round_up_dffe15 <= round_up_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe0 <= sign_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe1 <= sign_dffe0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe2 <= sign_dffe1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe3 <= sign_dffe2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe4 <= sign_dffe3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe5 <= sign_dffe4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe6 <= sign_dffe5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe7 <= sign_dffe6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe8 <= sign_dffe7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe9 <= sign_dffe8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe10 <= sign_dffe9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe11 <= sign_dffe10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe12 <= sign_dffe11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe13 <= sign_dffe12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe14 <= sign_dffe13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe15 <= sign_dffe14;
			END IF;
		END IF;
	END PROCESS;
	wire_sign_dffe_w_lg_q448w(0) <= sign_dffe15 AND wire_w_lg_distance_overflow447w(0);
	wire_sign_dffe_w_lg_q434w(0) <= NOT sign_dffe15;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN tbl1_compare_dffe11_4_pipes0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN tbl1_compare_dffe11_4_pipes0 <= tbl1_compare_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN tbl1_compare_dffe11_4_pipes1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN tbl1_compare_dffe11_4_pipes1 <= tbl1_compare_dffe11_4_pipes0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN tbl1_compare_dffe11_4_pipes2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN tbl1_compare_dffe11_4_pipes2 <= tbl1_compare_dffe11_4_pipes1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN tbl1_compare_dffe11_4_pipes3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN tbl1_compare_dffe11_4_pipes3 <= tbl1_compare_dffe11_4_pipes2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN tbl1_tbl2_prod_dffe12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN tbl1_tbl2_prod_dffe12 <= tbl1_tbl2_prod_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN tbl3_taylor_prod_dffe12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN tbl3_taylor_prod_dffe12 <= tbl3_taylor_prod_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_fixed_dffe_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_fixed_dffe_0 <= x_fixed;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_fixed_dffe_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_fixed_dffe_1 <= x_fixed_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_fixed_dffe_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_fixed_dffe_2 <= x_fixed_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_fixed_dffe_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_fixed_dffe_3 <= x_fixed_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_fixed_dffe_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_fixed_dffe_4 <= x_fixed_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN xf_pre_2_dffe10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN xf_pre_2_dffe10 <= xf_pre_2_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN xf_pre_dffe9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN xf_pre_dffe9 <= xf_pre_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN xi_exp_value_dffe4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN xi_exp_value_dffe4 <= xi_exp_value_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN xi_ln2_prod_dffe7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN xi_ln2_prod_dffe7 <= xi_ln2_prod_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN xi_prod_dffe3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN xi_prod_dffe3 <= xi_prod_wi;
			END IF;
		END IF;
	END PROCESS;
	wire_exp_minus_bias_dataa <= ( "0" & exp_w);
	wire_exp_minus_bias_datab <= ( "0" & exp_bias);
	exp_minus_bias :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => wire_exp_minus_bias_dataa,
		datab => wire_exp_minus_bias_datab,
		result => wire_exp_minus_bias_result
	  );
	wire_exp_value_add_bias_w_lg_w_result_range445w446w(0) <= NOT wire_exp_value_add_bias_w_result_range445w(0);
	wire_exp_value_add_bias_dataa <= ( "0" & exp_value_b4_bias_dffe_10);
	wire_exp_value_add_bias_datab <= ( "0" & exp_bias(7 DOWNTO 1) & wire_extra_ln2_dffe_5_w_lg_q157w);
	wire_exp_value_add_bias_w_result_range445w(0) <= wire_exp_value_add_bias_result(8);
	exp_value_add_bias :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_cin_to_bias_dataout,
		clken => clk_en,
		clock => clock,
		dataa => wire_exp_value_add_bias_dataa,
		datab => wire_exp_value_add_bias_datab,
		result => wire_exp_value_add_bias_result
	  );
	wire_exp_value_man_over_w_lg_w_lg_w_result_range435w436w437w(0) <= wire_exp_value_man_over_w_lg_w_result_range435w436w(0) AND wire_sign_dffe_w_lg_q434w(0);
	wire_exp_value_man_over_w_lg_w_result_range435w436w(0) <= NOT wire_exp_value_man_over_w_result_range435w(0);
	wire_exp_value_man_over_w_lg_w_lg_w_lg_w_result_range435w436w437w438w(0) <= wire_exp_value_man_over_w_lg_w_lg_w_result_range435w436w437w(0) OR sign_dffe15;
	wire_exp_value_man_over_datab <= ( "00000000" & man_overflow_wo);
	wire_exp_value_man_over_w_result_range435w(0) <= wire_exp_value_man_over_result(8);
	exp_value_man_over :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => wire_exp_value_add_bias_result,
		datab => wire_exp_value_man_over_datab,
		result => wire_exp_value_man_over_result
	  );
	wire_invert_exp_value_dataa <= (OTHERS => '0');
	wire_invert_exp_value_w_result_range130w <= wire_invert_exp_value_result(5 DOWNTO 0);
	invert_exp_value :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_invert_exp_value_dataa,
		datab => exp_value(7 DOWNTO 0),
		result => wire_invert_exp_value_result
	  );
	wire_man_round_datab <= ( "0000000000000000000000" & round_up_wo);
	man_round :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 23
	  )
	  PORT MAP ( 
		dataa => man_round_wo,
		datab => wire_man_round_datab,
		result => wire_man_round_result
	  );
	wire_one_minus_xf_dataa <= ( "1" & "000000000000000000000000000000");
	one_minus_xf :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 31
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_one_minus_xf_dataa,
		datab => wire_extra_ln2_muxa_dataout,
		result => wire_one_minus_xf_result
	  );
	wire_x_fixed_minus_xiln2_datab <= ( "0" & xi_ln2_prod_wo(45 DOWNTO 9));
	x_fixed_minus_xiln2 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 38
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => x_fixed_dffe_4,
		datab => wire_x_fixed_minus_xiln2_datab,
		result => wire_x_fixed_minus_xiln2_result
	  );
	wire_xf_minus_ln2_datab <= ( "00" & ln2_w(37 DOWNTO 9));
	xf_minus_ln2 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 31
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => xf_pre(30 DOWNTO 0),
		datab => wire_xf_minus_ln2_datab,
		result => wire_xf_minus_ln2_result
	  );
	wire_xi_add_one_datab <= "00000001";
	xi_add_one :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => xi_exp_value,
		datab => wire_xi_add_one_datab,
		result => wire_xi_add_one_result
	  );
	rbarrel_shift :  lpm_clshift
	  GENERIC MAP (
		LPM_PIPELINE => 2,
		LPM_SHIFTTYPE => "LOGICAL",
		LPM_WIDTH => 38,
		LPM_WIDTHDIST => 6
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		data => barrel_shifter_data,
		direction => exp_value_wo(8),
		distance => barrel_shifter_distance,
		result => wire_rbarrel_shift_result
	  );
	distance_overflow_comp :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		agb => wire_distance_overflow_comp_agb,
		dataa => wire_exp_value_to_compare_muxa_dataout,
		datab => distance_overflow_val_w
	  );
	tbl1_compare :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		ageb => wire_tbl1_compare_ageb,
		dataa => xf(28 DOWNTO 24),
		datab => addr_val_more_than_one
	  );
	underflow_compare :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		agb => wire_underflow_compare_agb,
		dataa => wire_exp_value_to_compare_muxa_dataout,
		datab => underflow_compare_val_w
	  );
	man_prod :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 31,
		LPM_WIDTHB => 31,
		LPM_WIDTHP => 62,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => tbl1_tbl2_prod_wo,
		datab => tbl3_taylor_prod_wo,
		result => wire_man_prod_result
	  );
	tbl1_tbl2_prod :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 32,
		LPM_WIDTHB => 32,
		LPM_WIDTHP => 64,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => table_one_out,
		datab => table_two_out,
		result => wire_tbl1_tbl2_prod_result
	  );
	wire_tbl3_taylor_prod_datab <= ( "1" & "000000000000000" & xf(13 DOWNTO 0));
	tbl3_taylor_prod :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 32,
		LPM_WIDTHB => 30,
		LPM_WIDTHP => 62,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => table_three_out,
		datab => wire_tbl3_taylor_prod_datab,
		result => wire_tbl3_taylor_prod_result
	  );
	xi_ln2_prod :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 2,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 8,
		LPM_WIDTHB => 38,
		LPM_WIDTHP => 46,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_exp_value_to_ln2a_dataout,
		datab => ln2_w,
		result => wire_xi_ln2_prod_result
	  );
	xi_prod :  lpm_mult
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 12,
		LPM_WIDTHB => 9,
		LPM_WIDTHP => 21,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		dataa => x_fixed(37 DOWNTO 26),
		datab => one_over_ln2_w,
		result => wire_xi_prod_result
	  );
	loop2 : FOR i IN 0 TO 31 GENERATE
		loop3 : FOR j IN 0 TO 31 GENERATE
			wire_table_one_data_2d(i, j) <= table_one_data(i*32+j);
		END GENERATE loop3;
	END GENERATE loop2;
	table_one :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 32,
		LPM_WIDTH => 32,
		LPM_WIDTHS => 5
	  )
	  PORT MAP ( 
		data => wire_table_one_data_2d,
		result => wire_table_one_result,
		sel => xf(28 DOWNTO 24)
	  );
	loop4 : FOR i IN 0 TO 31 GENERATE
		loop5 : FOR j IN 0 TO 20 GENERATE
			wire_table_three_data_2d(i, j) <= table_three_data(i*21+j);
		END GENERATE loop5;
	END GENERATE loop4;
	table_three :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 32,
		LPM_WIDTH => 21,
		LPM_WIDTHS => 5
	  )
	  PORT MAP ( 
		data => wire_table_three_data_2d,
		result => wire_table_three_result,
		sel => xf(18 DOWNTO 14)
	  );
	loop6 : FOR i IN 0 TO 31 GENERATE
		loop7 : FOR j IN 0 TO 25 GENERATE
			wire_table_two_data_2d(i, j) <= table_two_data(i*26+j);
		END GENERATE loop7;
	END GENERATE loop6;
	table_two :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 32,
		LPM_WIDTH => 26,
		LPM_WIDTHS => 5
	  )
	  PORT MAP ( 
		data => wire_table_two_data_2d,
		result => wire_table_two_result,
		sel => xf(23 DOWNTO 19)
	  );
	wire_cin_to_bias_dataout <= shifted_value;
	wire_exp_result_mux_prea_dataout <= exp_one WHEN wire_w_lg_w551w552w(0) = '1'  ELSE exp_result_w;
	loop8 : FOR i IN 0 TO 7 GENERATE 
		wire_exp_result_mux_prea_w_lg_dataout557w(i) <= wire_exp_result_mux_prea_dataout(i) AND wire_w_lg_w_lg_w_lg_underflow_w554w555w556w(0);
	END GENERATE loop8;
	wire_exp_value_b4_biasa_dataout <= exp_invert WHEN sign_dffe3 = '1'  ELSE xi_exp_value;
	wire_exp_value_selecta_dataout <= wire_invert_exp_value_result(5 DOWNTO 0) WHEN exp_value_wo(8) = '1'  ELSE exp_value_wo(5 DOWNTO 0);
	wire_exp_value_to_compare_muxa_dataout <= wire_invert_exp_value_result WHEN exp_value_wo(8) = '1'  ELSE exp_value_wo(7 DOWNTO 0);
	wire_exp_value_to_ln2a_dataout <= wire_xi_add_one_result WHEN sign_dffe4 = '1'  ELSE xi_exp_value_wo;
	wire_extra_ln2_muxa_dataout <= wire_xf_minus_ln2_result WHEN extra_ln2_dffe_0 = '1'  ELSE xf_pre_wo(30 DOWNTO 0);
	wire_man_result_muxa_dataout <= ( nan_w & "0000000000000000000000") WHEN wire_w_lg_w_lg_w_lg_w_lg_overflow_w536w537w538w539w(0) = '1'  ELSE wire_man_round_result;
	wire_xf_muxa_dataout <= wire_one_minus_xf_result WHEN sign_dffe10 = '1'  ELSE xf_pre_2_wo(30 DOWNTO 0);

 END RTL; --f_p_exp_altfp_exp_jmc
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY f_p_exp IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		data		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END f_p_exp;


ARCHITECTURE RTL OF f_p_exp IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT f_p_exp_altfp_exp_jmc
	PORT (
			clock	: IN STD_LOGIC ;
			data	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(31 DOWNTO 0);

	f_p_exp_altfp_exp_jmc_component : f_p_exp_altfp_exp_jmc
	PORT MAP (
		clock => clock,
		data => data,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altfp_exp"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "17"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "23"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: USED_PORT: data 0 0 32 0 INPUT NODEFVAL "data[31..0]"
-- Retrieval info: CONNECT: @data 0 0 32 0 data 0 0 32 0
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL f_p_exp.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL f_p_exp.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL f_p_exp.bsf TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL f_p_exp_inst.vhd TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL f_p_exp.inc TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL f_p_exp.cmp TRUE TRUE
-- Retrieval info: LIB_FILE: lpm

