f_p_exp_inst : f_p_exp PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		result	 => result_sig
	);
