f_p_inv_inst : f_p_inv PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		result	 => result_sig
	);
